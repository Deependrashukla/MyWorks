module notgate(a,c);
input a;
output c;
assign c=~a;
endmodule
